module or_gate_tb;
    reg a, b;
    wire y;

    //connect the OR gate
    or_gate uut (a, b, y);

    initial begin 
        $dumpfile("or_gate_results.vcd");
        $dumpvars(0, or_gate_tb);

        //truth table sequence 
        a=0; b=0; #10;
        a=0; b=1; #10;
        a=1; b=0; #10;
        a=1; b=1; #10;

        $display("OR gate tests complete");
        $finish;
    end
endmodule